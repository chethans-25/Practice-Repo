module fulladder()

endmodule